library verilog;
use verilog.vl_types.all;
entity test_xor is
end test_xor;
