library verilog;
use verilog.vl_types.all;
entity test_memory is
end test_memory;
