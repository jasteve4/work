library verilog;
use verilog.vl_types.all;
entity test_arbiter is
end test_arbiter;
